module beep_do (
	clk,
	o_do
);